class r_config extends uvm_object;
	`uvm_object_utils(r_config)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass
